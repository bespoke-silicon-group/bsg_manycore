
`include "bsg_manycore_defines.vh"

module bsg_manycore_link_ruche_to_sdr_west
 import bsg_noc_pkg::*;
 import bsg_manycore_pkg::*;
 #(parameter tieoff_east_not_west_p = 0
`include "bsg_manycore_link_ruche_to_sdr.vh"
endmodule

`BSG_ABSTRACT_MODULE(bsg_manycore_link_ruche_to_sdr_west)

