
`include "bsg_manycore_defines.svh"

module bsg_manycore_link_wh_to_sdr_se
`include "bsg_manycore_link_wh_to_sdr.svh"
endmodule

`BSG_ABSTRACT_MODULE(bsg_manycore_link_wh_to_sdr_se)

