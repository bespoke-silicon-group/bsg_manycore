module bsg_manycore_link_wh_to_sdr_nw
`include "bsg_manycore_link_wh_to_sdr.v"
endmodule