
`include "bsg_manycore_defines.vh"

module bsg_manycore_link_wh_to_sdr_ne
`include "bsg_manycore_link_wh_to_sdr.vh"
endmodule

`BSG_ABSTRACT_MODULE(bsg_manycore_link_wh_to_sdr_ne)

