module bsg_manycore_link_wh_to_sdr_se
`include "bsg_manycore_link_wh_to_sdr.v"
endmodule